`include "full_adder.sv"
`include "rca.sv"
module model (
    input [23:0] a,
    input [23:0] b,
    output logic [24:0] result
);

    

endmodule